module divb(clkin,clkout);
//input
input clkin;
//output
output reg clkout;
//reg&wire
reg [31:0]count;
wire [31:0]divn,divnh;

assign divn = 32'd3750000; //Frequency division ratio
assign divnh = divn>>1; //Half of divn

always@(posedge clkin)
begin
    if(count>=divn)
        count<=1;
    else
        count<=count+1;
end

always@(negedge clkin)
    clkout = (count<=divnh)?1:0;

endmodule